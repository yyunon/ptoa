-- Copyright 2018 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

-- This file was automatically generated by FletchGen. Modify this file
-- at your own risk.

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_misc.ALL;

LIBRARY work;
-- Fletcher
USE work.Interconnect_pkg.ALL;
USE work.Wrapper_pkg.ALL;

-- Ptoa
USE work.Ptoa.ALL;
ENTITY ptoa_wrapper IS
  GENERIC (
    BUS_ADDR_WIDTH : NATURAL;
    BUS_DATA_WIDTH : NATURAL;
    BUS_LEN_WIDTH : NATURAL;
    BUS_BURST_STEP_LEN : NATURAL;
    BUS_BURST_MAX_LEN : NATURAL;
    ---------------------------------------------------------------------------
    INDEX_WIDTH : NATURAL;
    ---------------------------------------------------------------------------
    NUM_ARROW_BUFFERS : NATURAL;
    NUM_REGS : NATURAL;
    REG_WIDTH : NATURAL;
    ---------------------------------------------------------------------------
    TAG_WIDTH : NATURAL
  );
  PORT (
    acc_reset : IN STD_LOGIC;
    bus_clk : IN STD_LOGIC;
    bus_reset : IN STD_LOGIC;
    acc_clk : IN STD_LOGIC;
    ---------------------------------------------------------------------------
    mst_rreq_valid : OUT STD_LOGIC;
    mst_rreq_ready : IN STD_LOGIC;
    mst_rreq_addr : OUT STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
    mst_rreq_len : OUT STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
    ---------------------------------------------------------------------------
    mst_rdat_valid : IN STD_LOGIC;
    mst_rdat_ready : OUT STD_LOGIC;
    mst_rdat_data : IN STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
    mst_rdat_last : IN STD_LOGIC;
    ---------------------------------------------------------------------------
    mst_wreq_valid : OUT STD_LOGIC;
    mst_wreq_len : OUT STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
    mst_wreq_last : OUT STD_LOGIC;
    mst_wreq_addr : OUT STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
    mst_wreq_ready : IN STD_LOGIC;
    ---------------------------------------------------------------------------
    mst_wdat_valid : OUT STD_LOGIC;
    mst_wdat_ready : IN STD_LOGIC;
    mst_wdat_data : OUT STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
    mst_wdat_strobe : OUT STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
    mst_wdat_last : OUT STD_LOGIC;
    ---------------------------------------------------------------------------
    regs_in : IN STD_LOGIC_VECTOR(NUM_REGS * REG_WIDTH - 1 DOWNTO 0);
    regs_out : OUT STD_LOGIC_VECTOR(NUM_REGS * REG_WIDTH - 1 DOWNTO 0);
    regs_out_en : OUT STD_LOGIC_VECTOR(NUM_REGS - 1 DOWNTO 0)
  );
END ptoa_wrapper;

ARCHITECTURE behv OF ptoa_wrapper IS
  ---------------------------------------
  -- Register offsets
  ---------------------------------------
  CONSTANT REG_CONTROL : NATURAL := 0;
  CONSTANT REG_STATUS : NATURAL := 1;

  --2 & 3 are return values
  --The following are schema-derived registers set by the fletcher runtime automatically, by queuing a recordbatch.
  -- See FLETCHER_REG_SCHEMA 
  CONSTANT REG_START_INDEX : NATURAL := 4;
  CONSTANT REG_END_INDEX : NATURAL := 5;
  CONSTANT REG_VAL_ADDR0 : NATURAL := 6;
  CONSTANT REG_VAL_ADDR1 : NATURAL := 7;
  --After the buffers needed for the record batch, the application code should set additional registers.
  --Coordinate these with REG_BASE in the application code.
  CONSTANT REG_NUM_VAL : NATURAL := 10;
  CONSTANT REG_PAGE_ADDR0 : NATURAL := 11;
  CONSTANT REG_PAGE_ADDR1 : NATURAL := 12;
  CONSTANT REG_MAX_SIZE0 : NATURAL := 13;
  CONSTANT REG_MAX_SIZE1 : NATURAL := 14;
  ---------------------------------------
  -- Fletcher UserCoreController signals
  ---------------------------------------
  SIGNAL uctrl_start : STD_LOGIC;
  SIGNAL uctrl_stop : STD_LOGIC;
  SIGNAL uctrl_reset : STD_LOGIC;
  SIGNAL uctrl_done : STD_LOGIC;

  ---------------------------------------
  -- Fletcher read/write arbiter signals
  ---------------------------------------
  SIGNAL bsv_rreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL bsv_rreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL bsv_rreq_ready : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL bsv_rreq_valid : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL bsv_rdat_valid : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL bsv_rdat_ready : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL bsv_rdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL bsv_rdat_last : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL bsv_wreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL bsv_wreq_last : STD_LOGIC;
  SIGNAL bsv_wreq_valid : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL bsv_wreq_ready : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL bsv_wreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);

  SIGNAL bsv_wrep_ready : STD_LOGIC;
  SIGNAL bsv_wrep_valid : STD_LOGIC;
  SIGNAL bsv_wrep_ok : STD_LOGIC;

  SIGNAL bsv_wdat_valid : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL bsv_wdat_last : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL bsv_wdat_strobe : STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL bsv_wdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL bsv_wdat_ready : STD_LOGIC_VECTOR(0 DOWNTO 0);

  -- ParquetReader reset
  SIGNAL pr_reset : STD_LOGIC;

  SIGNAL mst_wrep_valid : STD_LOGIC := '1';
  SIGNAL mst_wrep_ready : STD_LOGIC := '1';
  SIGNAL mst_wrep_ok : STD_LOGIC := '1';
BEGIN

  -- Only the status register needs to be written to
  regs_out_en <= (
    REG_CONTROL => '0',
    REG_STATUS => '1',
    REG_NUM_VAL => '0',
    REG_PAGE_ADDR0 => '0',
    REG_PAGE_ADDR1 => '0',
    REG_MAX_SIZE0 => '0',
    REG_MAX_SIZE1 => '0',
    REG_VAL_ADDR0 => '0',
    REG_VAL_ADDR1 => '0',
    OTHERS => '0');
  --  regs_out_en(REG_OFF_ADDR0)   <= '0';
  --  regs_out_en(REG_OFF_ADDR1)   <= '0';

  -- Reset the ParquetReader when the UserCoreController or the top level requests it
  pr_reset <= uctrl_reset OR bus_reset;

  -- Fletcher controller as a stand-in for future ptoa specific controller
  UserCoreController_inst : UserCoreController
  GENERIC MAP(
    REG_WIDTH => REG_WIDTH
  )
  PORT MAP(
    kcd_clk => acc_clk,
    kcd_reset => acc_reset,
    bcd_clk => bus_clk,
    bcd_reset => bus_reset,
    status => regs_out((REG_STATUS + 1) * REG_WIDTH - 1 DOWNTO REG_WIDTH * REG_STATUS),
    control => regs_in((REG_CONTROL + 1) * REG_WIDTH - 1 DOWNTO REG_WIDTH * REG_CONTROL),
    start => uctrl_start,
    stop => uctrl_stop,
    reset => uctrl_reset,
    idle => '0',
    busy => '0',
    done => uctrl_done
  );

  prim64_reader_inst : ParquetReader
  GENERIC MAP(
    BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    ---------------------------------------------------------------------------------
    INDEX_WIDTH => INDEX_WIDTH,
    ---------------------------------------------------------------------------------
    TAG_WIDTH => TAG_WIDTH,
    CFG => "prim(64;epc=8)",
    ENCODING => "DELTA",
    COMPRESSION_CODEC => "UNCOMPRESSED"
  )
  PORT MAP(
    clk => bus_clk,
    reset => pr_reset,
    bus_rreq_valid => bsv_rreq_valid(0),
    bus_rreq_ready => bsv_rreq_ready(0),
    bus_rreq_addr => bsv_rreq_addr,
    bus_rreq_len => bsv_rreq_len,
    bus_rdat_valid => bsv_rdat_valid(0),
    bus_rdat_ready => bsv_rdat_ready(0),
    bus_rdat_data => bsv_rdat_data,
    bus_rdat_last => bsv_rdat_last(0),
    bus_wreq_valid => bsv_wreq_valid(0),
    bus_wreq_len => bsv_wreq_len,
    bus_wreq_last => bsv_wreq_last,
    bus_wreq_addr => bsv_wreq_addr,
    bus_wreq_ready => bsv_wreq_ready(0),
    bus_wrep_valid => bsv_wrep_valid,
    bus_wrep_ready => bsv_wrep_ready,
    bus_wrep_ok => bsv_wrep_ok,
    bus_wdat_valid => bsv_wdat_valid(0),
    bus_wdat_ready => bsv_wdat_ready(0),
    bus_wdat_data => bsv_wdat_data,
    bus_wdat_strobe => bsv_wdat_strobe,
    bus_wdat_last => bsv_wdat_last(0),
    base_pages_ptr => regs_in((REG_PAGE_ADDR1 + 1) * REG_WIDTH - 1 DOWNTO REG_WIDTH * REG_PAGE_ADDR0),
    max_data_size => regs_in((REG_MAX_SIZE1 + 1) * REG_WIDTH - 1 DOWNTO REG_WIDTH * REG_MAX_SIZE0),
    total_num_values => regs_in((REG_NUM_VAL + 1) * REG_WIDTH - 1 DOWNTO REG_WIDTH * REG_NUM_VAL),
    values_buffer_addr => regs_in((REG_VAL_ADDR1 + 1) * REG_WIDTH - 1 DOWNTO REG_WIDTH * REG_VAL_ADDR0),
    offsets_buffer_addr => (OTHERS => '0'),
    start => uctrl_start,
    stop => uctrl_stop,
    done => uctrl_done
  );

  -- Fletcher BusWriteArbiter
  BusWriteArbiterVec_inst : BusWriteArbiterVec
  GENERIC MAP(
    BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    NUM_SLAVE_PORTS => 1,
    MAX_OUTSTANDING => 16
  )
  PORT MAP(
    bcd_clk => bus_clk,
    bcd_reset => bus_reset,
    bsv_wdat_valid => bsv_wdat_valid,
    bsv_wdat_ready => bsv_wdat_ready,
    bsv_wdat_data => bsv_wdat_data,
    bsv_wdat_strobe => bsv_wdat_strobe,
    bsv_wdat_last => bsv_wdat_last,
    bsv_wrep_valid(0) => bsv_wrep_valid,
    bsv_wrep_ready(0) => bsv_wrep_ready,
    bsv_wrep_ok(0) => bsv_wrep_ok,
    bsv_wreq_valid => bsv_wreq_valid,
    bsv_wreq_ready => bsv_wreq_ready,
    bsv_wreq_addr => bsv_wreq_addr,
    bsv_wreq_len => bsv_wreq_len,
    bsv_wreq_last(0) => bsv_wreq_last,
    mst_wreq_valid => mst_wreq_valid,
    mst_wreq_ready => mst_wreq_ready,
    mst_wreq_addr => mst_wreq_addr,
    mst_wreq_len => mst_wreq_len,
    mst_wreq_last => mst_wreq_last,
    mst_wdat_valid => mst_wdat_valid,
    mst_wdat_ready => mst_wdat_ready,
    mst_wdat_data => mst_wdat_data,
    mst_wdat_strobe => mst_wdat_strobe,
    mst_wdat_last => mst_wdat_last,
    mst_wrep_valid => mst_wrep_valid,
    mst_wrep_ready => mst_wrep_ready,
    mst_wrep_ok => mst_wrep_ok
  );

  -- Fletcher BusReadArbiter
  BusReadArbiterVec_inst : BusReadArbiterVec
  GENERIC MAP(
    BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    NUM_SLAVE_PORTS => 1,
    MAX_OUTSTANDING => 16
  )
  PORT MAP(
    bcd_clk => bus_clk,
    bcd_reset => bus_reset,
    bsv_rreq_valid => bsv_rreq_valid,
    bsv_rreq_ready => bsv_rreq_ready,
    bsv_rreq_addr => bsv_rreq_addr,
    bsv_rreq_len => bsv_rreq_len,
    bsv_rdat_valid => bsv_rdat_valid,
    bsv_rdat_ready => bsv_rdat_ready,
    bsv_rdat_data => bsv_rdat_data,
    bsv_rdat_last => bsv_rdat_last,
    mst_rreq_valid => mst_rreq_valid,
    mst_rreq_ready => mst_rreq_ready,
    mst_rreq_addr => mst_rreq_addr,
    mst_rreq_len => mst_rreq_len,
    mst_rdat_valid => mst_rdat_valid,
    mst_rdat_ready => mst_rdat_ready,
    mst_rdat_data => mst_rdat_data,
    mst_rdat_last => mst_rdat_last
  );

END ARCHITECTURE;